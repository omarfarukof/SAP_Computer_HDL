module ram (
    input R_W,
    input EnOut,
    input [3:0] Addr,
    input [7:0] DataIn,
    output [7:0] DataOut
);
    reg [7:0] reg [15:0];

    // ... ... ... 
    
endmodule